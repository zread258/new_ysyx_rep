module ysyx_23060184_IFU (
    input                           clk,
    input                           rstn,
    input [`DATA_WIDTH - 1:0]       NPC,
    input                           Evalid,
    output reg                      Eready,
    output reg                      Ivalid,
    output reg [`DATA_WIDTH - 1:0]  PC
);

endmodule